<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-29.5,-20.9192,309.454,-188.458</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>13.5,-2.5</position>
<gparam>LABEL_TEXT Asynchronous(RIPPLE) Counters</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>18.5,-6.5</position>
<gparam>LABEL_TEXT 1. 3 bit Up Counter(+ve edge triggering) : </gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>BE_JKFF_LOW</type>
<position>7.5,-19.5</position>
<input>
<ID>J</ID>1 </input>
<input>
<ID>K</ID>1 </input>
<output>
<ID>Q</ID>5 </output>
<input>
<ID>clock</ID>2 </input>
<output>
<ID>nQ</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>BE_JKFF_LOW</type>
<position>19.5,-19.5</position>
<input>
<ID>J</ID>1 </input>
<input>
<ID>K</ID>1 </input>
<output>
<ID>Q</ID>6 </output>
<input>
<ID>clock</ID>3 </input>
<output>
<ID>nQ</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>BE_JKFF_LOW</type>
<position>30.5,-19.5</position>
<input>
<ID>J</ID>1 </input>
<input>
<ID>K</ID>1 </input>
<output>
<ID>Q</ID>7 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-9,-13.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>BB_CLOCK</type>
<position>-9.5,-19.5</position>
<output>
<ID>CLK</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>16</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>43,-20</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>11.5,-11</position>
<input>
<ID>N_in2</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>23.5,-11</position>
<input>
<ID>N_in2</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>34,-11</position>
<input>
<ID>N_in2</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>19,-30</position>
<gparam>LABEL_TEXT 2. 3 bit Down Counter(+ve edge triggering) :</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>BE_JKFF_LOW</type>
<position>8,-44.5</position>
<input>
<ID>J</ID>8 </input>
<input>
<ID>K</ID>8 </input>
<output>
<ID>Q</ID>10 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>BE_JKFF_LOW</type>
<position>20,-44.5</position>
<input>
<ID>J</ID>8 </input>
<input>
<ID>K</ID>8 </input>
<output>
<ID>Q</ID>11 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>30</ID>
<type>BE_JKFF_LOW</type>
<position>33,-44.5</position>
<input>
<ID>J</ID>8 </input>
<input>
<ID>K</ID>8 </input>
<output>
<ID>Q</ID>15 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-6.5,-40.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>13.5,-35.5</position>
<input>
<ID>N_in2</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>24.5,-35.5</position>
<input>
<ID>N_in2</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>38,-35.5</position>
<input>
<ID>N_in2</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>43.5,-45</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>15 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>42</ID>
<type>BB_CLOCK</type>
<position>-6.5,-44.5</position>
<output>
<ID>CLK</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>17.5,-56</position>
<gparam>LABEL_TEXT 3. 4 bit up Counter(-ve edge Triggering) : </gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>BE_JKFF_LOW_NT</type>
<position>8,-70</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>17 </input>
<output>
<ID>Q</ID>22 </output>
<input>
<ID>clock</ID>18 </input>
<output>
<ID>nQ</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>BE_JKFF_LOW_NT</type>
<position>21,-70</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>17 </input>
<output>
<ID>Q</ID>23 </output>
<input>
<ID>clock</ID>19 </input>
<output>
<ID>nQ</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>50</ID>
<type>BE_JKFF_LOW_NT</type>
<position>34,-70</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>17 </input>
<output>
<ID>Q</ID>24 </output>
<input>
<ID>clock</ID>20 </input>
<output>
<ID>nQ</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>-6,-64.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>54</ID>
<type>BB_CLOCK</type>
<position>-7.5,-70</position>
<output>
<ID>CLK</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>56</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>62.5,-71</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<input>
<ID>IN_2</ID>23 </input>
<input>
<ID>IN_3</ID>22 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>-1,-78</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>60</ID>
<type>DE_TO</type>
<position>13,-78.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>62</ID>
<type>DE_TO</type>
<position>26,-78.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>64</ID>
<type>DE_TO</type>
<position>39,-78.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>66</ID>
<type>BE_JKFF_LOW_NT</type>
<position>46,-70</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>17 </input>
<output>
<ID>Q</ID>25 </output>
<input>
<ID>clock</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>68</ID>
<type>DE_TO</type>
<position>51,-79</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>13,-74.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>GA_LED</type>
<position>27,-75</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>40.5,-75.5</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>51.5,-75</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>21.5,-92</position>
<gparam>LABEL_TEXT 4. 4 Bit Up Down Counter(+ve edge triggering) :</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>BE_JKFF_LOW</type>
<position>3.5,-113.5</position>
<input>
<ID>J</ID>46 </input>
<input>
<ID>K</ID>46 </input>
<output>
<ID>Q</ID>38 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>111</ID>
<type>BE_JKFF_LOW</type>
<position>16.5,-113.5</position>
<input>
<ID>J</ID>46 </input>
<input>
<ID>K</ID>46 </input>
<output>
<ID>Q</ID>39 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>112</ID>
<type>BE_JKFF_LOW</type>
<position>29,-113.5</position>
<input>
<ID>J</ID>46 </input>
<input>
<ID>K</ID>46 </input>
<output>
<ID>Q</ID>40 </output>
<input>
<ID>clock</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_TOGGLE</type>
<position>-4.5,-102</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_TOGGLE</type>
<position>-6.5,-120</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>115</ID>
<type>BB_CLOCK</type>
<position>-10,-113.5</position>
<output>
<ID>CLK</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>9,-122</position>
<input>
<ID>N_in3</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>GA_LED</type>
<position>22.5,-122</position>
<input>
<ID>N_in3</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>36,-122</position>
<input>
<ID>N_in3</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>BE_JKFF_LOW</type>
<position>41.5,-113.5</position>
<input>
<ID>J</ID>46 </input>
<input>
<ID>K</ID>46 </input>
<output>
<ID>Q</ID>41 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>48,-122</position>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AO_XNOR2</type>
<position>10,-106</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AO_XNOR2</type>
<position>22.5,-106</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AO_XNOR2</type>
<position>35,-106</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>53.5,-113.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>41 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 14</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-21.5,-1,-13.5</points>
<intersection>-21.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-21.5,4.5,-21.5</points>
<connection>
<GID>6</GID>
<name>K</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7,-13.5,25.5,-13.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection>
<intersection>4.5 8</intersection>
<intersection>14.5 7</intersection>
<intersection>16.5 14</intersection>
<intersection>25.5 13</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>14.5,-21.5,14.5,-13.5</points>
<intersection>-21.5 10</intersection>
<intersection>-13.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>4.5,-17.5,4.5,-13.5</points>
<connection>
<GID>6</GID>
<name>J</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>14.5,-21.5,16.5,-21.5</points>
<connection>
<GID>8</GID>
<name>K</name></connection>
<intersection>14.5 7</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>25.5,-21.5,25.5,-13.5</points>
<intersection>-21.5 16</intersection>
<intersection>-17.5 17</intersection>
<intersection>-13.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>16.5,-17.5,16.5,-13.5</points>
<connection>
<GID>8</GID>
<name>J</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>25.5,-21.5,27.5,-21.5</points>
<connection>
<GID>10</GID>
<name>K</name></connection>
<intersection>25.5 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>25.5,-17.5,27.5,-17.5</points>
<connection>
<GID>10</GID>
<name>J</name></connection>
<intersection>25.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-19.5,4.5,-19.5</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<connection>
<GID>14</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-21.5,13.5,-19.5</points>
<intersection>-21.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-19.5,16.5,-19.5</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-21.5,13.5,-21.5</points>
<connection>
<GID>6</GID>
<name>nQ</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-21.5,25,-19.5</points>
<intersection>-21.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-19.5,27.5,-19.5</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-21.5,25,-21.5</points>
<connection>
<GID>8</GID>
<name>nQ</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-26,11.5,-12</points>
<connection>
<GID>18</GID>
<name>N_in2</name></connection>
<intersection>-26 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-17.5,11.5,-17.5</points>
<connection>
<GID>6</GID>
<name>Q</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-26,40,-26</points>
<intersection>11.5 0</intersection>
<intersection>40 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-26,40,-21</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-26 2</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-24.5,23.5,-12</points>
<connection>
<GID>20</GID>
<name>N_in2</name></connection>
<intersection>-24.5 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-17.5,23.5,-17.5</points>
<connection>
<GID>8</GID>
<name>Q</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-24.5,38,-24.5</points>
<intersection>23.5 0</intersection>
<intersection>38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-24.5,38,-20</points>
<intersection>-24.5 2</intersection>
<intersection>-20 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38,-20,40,-20</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-19,34,-12</points>
<connection>
<GID>22</GID>
<name>N_in2</name></connection>
<intersection>-19 4</intersection>
<intersection>-17.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-17.5,34,-17.5</points>
<connection>
<GID>10</GID>
<name>Q</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>34,-19,40,-19</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-46.5,0,-40.5</points>
<intersection>-46.5 4</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-40.5,30,-40.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>0 0</intersection>
<intersection>5 7</intersection>
<intersection>17 6</intersection>
<intersection>30 12</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>0,-46.5,5,-46.5</points>
<connection>
<GID>26</GID>
<name>K</name></connection>
<intersection>0 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>17,-46.5,17,-40.5</points>
<connection>
<GID>28</GID>
<name>K</name></connection>
<connection>
<GID>28</GID>
<name>J</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>5,-42.5,5,-40.5</points>
<connection>
<GID>26</GID>
<name>J</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>30,-46.5,30,-40.5</points>
<connection>
<GID>30</GID>
<name>K</name></connection>
<connection>
<GID>30</GID>
<name>J</name></connection>
<intersection>-40.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-44.5,5,-44.5</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<connection>
<GID>42</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-49.5,12,-42.5</points>
<intersection>-49.5 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-49.5,40.5,-49.5</points>
<intersection>12 0</intersection>
<intersection>14 4</intersection>
<intersection>40.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-42.5,13.5,-42.5</points>
<connection>
<GID>26</GID>
<name>Q</name></connection>
<intersection>12 0</intersection>
<intersection>13.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40.5,-49.5,40.5,-46</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>14,-49.5,14,-44.5</points>
<intersection>-49.5 1</intersection>
<intersection>-44.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>13.5,-42.5,13.5,-36.5</points>
<connection>
<GID>34</GID>
<name>N_in2</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>14,-44.5,17,-44.5</points>
<connection>
<GID>28</GID>
<name>clock</name></connection>
<intersection>14 4</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-48.5,26.5,-42.5</points>
<intersection>-48.5 1</intersection>
<intersection>-44.5 9</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-48.5,39,-48.5</points>
<intersection>26.5 0</intersection>
<intersection>39 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-42.5,26.5,-42.5</points>
<connection>
<GID>28</GID>
<name>Q</name></connection>
<intersection>24.5 5</intersection>
<intersection>26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39,-48.5,39,-45</points>
<intersection>-48.5 1</intersection>
<intersection>-45 7</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>24.5,-42.5,24.5,-36.5</points>
<connection>
<GID>36</GID>
<name>N_in2</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>39,-45,40.5,-45</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>39 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>26.5,-44.5,30,-44.5</points>
<connection>
<GID>30</GID>
<name>clock</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-44,38,-36.5</points>
<connection>
<GID>38</GID>
<name>N_in2</name></connection>
<intersection>-44 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-44,40.5,-44</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-42.5,38,-42.5</points>
<connection>
<GID>30</GID>
<name>Q</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-64.5,42.5,-64.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>3.5 4</intersection>
<intersection>18 9</intersection>
<intersection>31 13</intersection>
<intersection>42.5 17</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>3.5,-72,3.5,-64.5</points>
<intersection>-72 6</intersection>
<intersection>-68 15</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>3.5,-72,5,-72</points>
<connection>
<GID>46</GID>
<name>K</name></connection>
<intersection>3.5 4</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>18,-72,18,-64.5</points>
<connection>
<GID>48</GID>
<name>K</name></connection>
<connection>
<GID>48</GID>
<name>J</name></connection>
<intersection>-64.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>31,-72,31,-64.5</points>
<connection>
<GID>50</GID>
<name>K</name></connection>
<connection>
<GID>50</GID>
<name>J</name></connection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>3.5,-68,5,-68</points>
<connection>
<GID>46</GID>
<name>J</name></connection>
<intersection>3.5 4</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>42.5,-72,42.5,-64.5</points>
<intersection>-72 19</intersection>
<intersection>-68 20</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>42.5,-72,43,-72</points>
<connection>
<GID>66</GID>
<name>K</name></connection>
<intersection>42.5 17</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>42.5,-68,43,-68</points>
<connection>
<GID>66</GID>
<name>J</name></connection>
<intersection>42.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,-70,5,-70</points>
<connection>
<GID>46</GID>
<name>clock</name></connection>
<connection>
<GID>54</GID>
<name>CLK</name></connection>
<intersection>-3 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-3,-78,-3,-70</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-70 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-72,14.5,-70</points>
<intersection>-72 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-70,18,-70</points>
<connection>
<GID>48</GID>
<name>clock</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-72,14.5,-72</points>
<connection>
<GID>46</GID>
<name>nQ</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-72,27.5,-70</points>
<intersection>-72 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-70,31,-70</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-72,27.5,-72</points>
<connection>
<GID>48</GID>
<name>nQ</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-72,40,-70</points>
<intersection>-72 1</intersection>
<intersection>-70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-72,40,-72</points>
<connection>
<GID>50</GID>
<name>nQ</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-70,43,-70</points>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-84.5,11,-68</points>
<connection>
<GID>46</GID>
<name>Q</name></connection>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-84.5 4</intersection>
<intersection>-74.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>11,-84.5,55.5,-84.5</points>
<intersection>11 0</intersection>
<intersection>55.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>55.5,-84.5,55.5,-69</points>
<intersection>-84.5 4</intersection>
<intersection>-69 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>11,-74.5,12,-74.5</points>
<connection>
<GID>70</GID>
<name>N_in0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>55.5,-69,59.5,-69</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>55.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-86,24,-68</points>
<connection>
<GID>48</GID>
<name>Q</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-86 1</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-86,56.5,-86</points>
<intersection>24 0</intersection>
<intersection>56.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>56.5,-86,56.5,-70</points>
<intersection>-86 1</intersection>
<intersection>-70 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24,-75,26,-75</points>
<connection>
<GID>72</GID>
<name>N_in0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>56.5,-70,59.5,-70</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>56.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-87.5,37,-68</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>Q</name></connection>
<intersection>-87.5 4</intersection>
<intersection>-75.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-87.5,57.5,-87.5</points>
<intersection>37 0</intersection>
<intersection>57.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>57.5,-87.5,57.5,-71</points>
<intersection>-87.5 4</intersection>
<intersection>-71 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>37,-75.5,39.5,-75.5</points>
<connection>
<GID>74</GID>
<name>N_in0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>57.5,-71,59.5,-71</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>57.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-88.5,49,-68</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<connection>
<GID>66</GID>
<name>Q</name></connection>
<intersection>-88.5 1</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-88.5,58.5,-88.5</points>
<intersection>49 0</intersection>
<intersection>58.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>58.5,-88.5,58.5,-72</points>
<intersection>-88.5 1</intersection>
<intersection>-72 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>49,-75,50.5,-75</points>
<connection>
<GID>76</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>58.5,-72,59.5,-72</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>58.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-113.5,0.5,-113.5</points>
<connection>
<GID>115</GID>
<name>CLK</name></connection>
<connection>
<GID>110</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-121,9,-111.5</points>
<connection>
<GID>116</GID>
<name>N_in3</name></connection>
<intersection>-120.5 4</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-111.5,9,-111.5</points>
<connection>
<GID>110</GID>
<name>Q</name></connection>
<intersection>7 2</intersection>
<intersection>9 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>7,-111.5,7,-107</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>9,-120.5,50,-120.5</points>
<intersection>9 0</intersection>
<intersection>50 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>50,-120.5,50,-114.5</points>
<intersection>-120.5 4</intersection>
<intersection>-114.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>50,-114.5,50.5,-114.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>50 5</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-121,22.5,-111.5</points>
<connection>
<GID>117</GID>
<name>N_in3</name></connection>
<intersection>-120 3</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-111.5,22.5,-111.5</points>
<connection>
<GID>111</GID>
<name>Q</name></connection>
<intersection>19.5 2</intersection>
<intersection>22.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>19.5,-111.5,19.5,-107</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-120,49.5,-120</points>
<intersection>22.5 0</intersection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-120,49.5,-113.5</points>
<intersection>-120 3</intersection>
<intersection>-113.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>49.5,-113.5,50.5,-113.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>49.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-121,36,-111.5</points>
<connection>
<GID>118</GID>
<name>N_in3</name></connection>
<intersection>-119.5 3</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-111.5,36,-111.5</points>
<connection>
<GID>112</GID>
<name>Q</name></connection>
<intersection>32 2</intersection>
<intersection>36 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>32,-111.5,32,-107</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>36,-119.5,49,-119.5</points>
<intersection>36 0</intersection>
<intersection>49 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49,-119.5,49,-112.5</points>
<intersection>-119.5 3</intersection>
<intersection>-112.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>49,-112.5,50.5,-112.5</points>
<connection>
<GID>124</GID>
<name>IN_2</name></connection>
<intersection>49 4</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-121,48,-111.5</points>
<connection>
<GID>120</GID>
<name>N_in3</name></connection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-111.5,50.5,-111.5</points>
<connection>
<GID>124</GID>
<name>IN_3</name></connection>
<connection>
<GID>119</GID>
<name>Q</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-102,32,-102</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>7 7</intersection>
<intersection>19.5 6</intersection>
<intersection>32 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>32,-105,32,-102</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>-102 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>19.5,-105,19.5,-102</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-102 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>7,-105,7,-102</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>-102 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-113.5,13,-106</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-113.5,13.5,-113.5</points>
<connection>
<GID>111</GID>
<name>clock</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-113.5,25.5,-106</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-113.5,26,-113.5</points>
<connection>
<GID>112</GID>
<name>clock</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-113.5,38,-106</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-113.5,38.5,-113.5</points>
<connection>
<GID>119</GID>
<name>clock</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-120,-1.5,-115.5</points>
<intersection>-120 1</intersection>
<intersection>-115.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-120,37,-120</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection>
<intersection>0.5 7</intersection>
<intersection>12.5 6</intersection>
<intersection>25 11</intersection>
<intersection>37 17</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1.5,-115.5,0.5,-115.5</points>
<connection>
<GID>110</GID>
<name>K</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>12.5,-120,12.5,-111.5</points>
<intersection>-120 1</intersection>
<intersection>-115.5 9</intersection>
<intersection>-111.5 13</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>0.5,-120,0.5,-111.5</points>
<connection>
<GID>110</GID>
<name>J</name></connection>
<intersection>-120 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>12.5,-115.5,13.5,-115.5</points>
<connection>
<GID>111</GID>
<name>K</name></connection>
<intersection>12.5 6</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>25,-120,25,-111.5</points>
<intersection>-120 1</intersection>
<intersection>-115.5 15</intersection>
<intersection>-111.5 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>12.5,-111.5,13.5,-111.5</points>
<connection>
<GID>111</GID>
<name>J</name></connection>
<intersection>12.5 6</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>25,-115.5,26,-115.5</points>
<connection>
<GID>112</GID>
<name>K</name></connection>
<intersection>25 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>37,-120,37,-111.5</points>
<intersection>-120 1</intersection>
<intersection>-115.5 21</intersection>
<intersection>-111.5 20</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>25,-111.5,26,-111.5</points>
<connection>
<GID>112</GID>
<name>J</name></connection>
<intersection>25 11</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>37,-111.5,38.5,-111.5</points>
<connection>
<GID>119</GID>
<name>J</name></connection>
<intersection>37 17</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>37,-115.5,38.5,-115.5</points>
<connection>
<GID>119</GID>
<name>K</name></connection>
<intersection>37 17</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>15.3,26.6356,269.515,-99.0183</PageViewport>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>45.5,-0.5</position>
<gparam>LABEL_TEXT Synchronous Counter </gparam>
<gparam>TEXT_HEIGHT 1.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>41.5,-5.5</position>
<gparam>LABEL_TEXT 3 Bit Up Counter</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>BE_JKFF_LOW</type>
<position>34,-25</position>
<input>
<ID>J</ID>48 </input>
<input>
<ID>K</ID>48 </input>
<output>
<ID>Q</ID>49 </output>
<input>
<ID>clock</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>132</ID>
<type>BE_JKFF_LOW</type>
<position>49,-25</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>50 </output>
<input>
<ID>clock</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>134</ID>
<type>BE_JKFF_LOW</type>
<position>63.5,-25</position>
<input>
<ID>J</ID>51 </input>
<output>
<ID>Q</ID>52 </output>
<input>
<ID>clock</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_AND2</type>
<position>56,-17</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>39.5,-33</position>
<input>
<ID>N_in3</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>GA_LED</type>
<position>54,-33</position>
<input>
<ID>N_in3</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>GA_LED</type>
<position>68.5,-33</position>
<input>
<ID>N_in3</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>BB_CLOCK</type>
<position>21.5,-30.5</position>
<output>
<ID>CLK</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>150</ID>
<type>EE_VDD</type>
<position>26.5,-18</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-30.5,60.5,-30.5</points>
<connection>
<GID>148</GID>
<name>CLK</name></connection>
<intersection>29.5 5</intersection>
<intersection>46 4</intersection>
<intersection>60.5 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46,-30.5,46,-25</points>
<connection>
<GID>132</GID>
<name>clock</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>29.5,-30.5,29.5,-25</points>
<intersection>-30.5 1</intersection>
<intersection>-25 8</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>60.5,-30.5,60.5,-25</points>
<connection>
<GID>134</GID>
<name>clock</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>29.5,-25,31,-25</points>
<connection>
<GID>130</GID>
<name>clock</name></connection>
<intersection>29.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-27,26.5,-19</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>-27 4</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-23,31,-23</points>
<connection>
<GID>130</GID>
<name>J</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-27,31,-27</points>
<connection>
<GID>130</GID>
<name>K</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-23,46,-23</points>
<connection>
<GID>132</GID>
<name>J</name></connection>
<connection>
<GID>130</GID>
<name>Q</name></connection>
<intersection>39.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,-32,39.5,-16</points>
<connection>
<GID>142</GID>
<name>N_in3</name></connection>
<intersection>-27 4</intersection>
<intersection>-23 1</intersection>
<intersection>-16 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>39.5,-27,46,-27</points>
<connection>
<GID>132</GID>
<name>K</name></connection>
<intersection>39.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>39.5,-16,53,-16</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>39.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-32,54,-23</points>
<connection>
<GID>144</GID>
<name>N_in3</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-23,54,-23</points>
<connection>
<GID>132</GID>
<name>Q</name></connection>
<intersection>52 2</intersection>
<intersection>54 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>52,-23,52,-18</points>
<intersection>-23 1</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-18,53,-18</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>52 2</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-23,59.5,-17</points>
<intersection>-23 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-23,60.5,-23</points>
<connection>
<GID>134</GID>
<name>J</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-17,59.5,-17</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-32,68.5,-23</points>
<connection>
<GID>146</GID>
<name>N_in3</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-23,68.5,-23</points>
<connection>
<GID>134</GID>
<name>Q</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>15.3,26.6356,269.515,-99.0183</PageViewport>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>54,-2.5</position>
<gparam>LABEL_TEXT SISO Shift Right</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>BB_CLOCK</type>
<position>25,-30.5</position>
<output>
<ID>CLK</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>170</ID>
<type>GA_LED</type>
<position>43.5,-15</position>
<input>
<ID>N_in2</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>GA_LED</type>
<position>55.5,-15</position>
<input>
<ID>N_in2</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>GA_LED</type>
<position>67,-15</position>
<input>
<ID>N_in2</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>GA_LED</type>
<position>77,-15</position>
<input>
<ID>N_in2</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AE_DFF_LOW</type>
<position>39.5,-23</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>61 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>184</ID>
<type>AE_DFF_LOW</type>
<position>51.5,-22.5</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>63 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_DFF_LOW</type>
<position>62,-22.5</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>188</ID>
<type>AE_DFF_LOW</type>
<position>73,-22.5</position>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>190</ID>
<type>BB_CLOCK</type>
<position>25.5,-21.5</position>
<output>
<ID>CLK</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 7</lparam></gate>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-21,43.5,-16</points>
<connection>
<GID>170</GID>
<name>N_in2</name></connection>
<intersection>-21 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-21,43.5,-21</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-20.5,48.5,-20.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-30.5,70,-30.5</points>
<connection>
<GID>168</GID>
<name>CLK</name></connection>
<intersection>36.5 8</intersection>
<intersection>48.5 3</intersection>
<intersection>59 7</intersection>
<intersection>70 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-30.5,48.5,-23.5</points>
<connection>
<GID>184</GID>
<name>clock</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>70,-30.5,70,-23.5</points>
<connection>
<GID>188</GID>
<name>clock</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>59,-30.5,59,-23.5</points>
<connection>
<GID>186</GID>
<name>clock</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>36.5,-30.5,36.5,-24</points>
<connection>
<GID>182</GID>
<name>clock</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-20.5,59,-20.5</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>55.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55.5,-20.5,55.5,-16</points>
<connection>
<GID>172</GID>
<name>N_in2</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-20.5,67,-16</points>
<connection>
<GID>174</GID>
<name>N_in2</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-20.5,70,-20.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-20.5,77,-16</points>
<connection>
<GID>176</GID>
<name>N_in2</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-20.5,77,-20.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-21.5,33,-21</points>
<intersection>-21.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-21,36.5,-21</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-21.5,33,-21.5</points>
<connection>
<GID>190</GID>
<name>CLK</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>9.3,31.1356,263.515,-94.5183</PageViewport>
<gate>
<ID>194</ID>
<type>AE_DFF_LOW</type>
<position>38,-24</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>81 </output>
<input>
<ID>clock</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_DFF_LOW</type>
<position>50,-24</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>82 </output>
<input>
<ID>clock</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>198</ID>
<type>AE_DFF_LOW</type>
<position>62.5,-24</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>83 </output>
<input>
<ID>clock</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_DFF_LOW</type>
<position>74,-24</position>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>84 </output>
<input>
<ID>clock</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_TOGGLE</type>
<position>26,-6.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>204</ID>
<type>BB_CLOCK</type>
<position>25.5,-30</position>
<output>
<ID>CLK</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_AND2</type>
<position>29,-12.5</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_AND2</type>
<position>33.5,-12.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_OR2</type>
<position>31.5,-19</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>42,-12.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_AND2</type>
<position>46.5,-12.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_OR2</type>
<position>44.5,-19</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>54,-12.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_AND2</type>
<position>58.5,-12.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AE_OR2</type>
<position>56.5,-19</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_AND2</type>
<position>66,-12.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>70.5,-12.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AE_OR2</type>
<position>68.5,-19</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_INVERTER</type>
<position>36.5,-3</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>223</ID>
<type>GA_LED</type>
<position>42,-34.5</position>
<input>
<ID>N_in3</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>GA_LED</type>
<position>54,-34.5</position>
<input>
<ID>N_in3</ID>82 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>GA_LED</type>
<position>66,-35</position>
<input>
<ID>N_in3</ID>83 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>229</ID>
<type>GA_LED</type>
<position>79,-35.5</position>
<input>
<ID>N_in3</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_TOGGLE</type>
<position>30,-7.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_TOGGLE</type>
<position>69.5,-7.5</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>52,-31.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID q2</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>64,-32</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID q3</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>77,-32.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID q4</lparam></gate>
<gate>
<ID>243</ID>
<type>DE_TO</type>
<position>32.5,-7.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID q2</lparam></gate>
<gate>
<ID>244</ID>
<type>DE_TO</type>
<position>45.5,-7.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID q3</lparam></gate>
<gate>
<ID>245</ID>
<type>DE_TO</type>
<position>57.5,-7.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID q4</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>48,1</position>
<gparam>LABEL_TEXT Bidirectional Registor : </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-30,71,-30</points>
<connection>
<GID>204</GID>
<name>CLK</name></connection>
<intersection>35 8</intersection>
<intersection>47 3</intersection>
<intersection>59.5 7</intersection>
<intersection>71 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47,-30,47,-25</points>
<connection>
<GID>196</GID>
<name>clock</name></connection>
<intersection>-30 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>71,-30,71,-25</points>
<connection>
<GID>200</GID>
<name>clock</name></connection>
<intersection>-30 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>59.5,-30,59.5,-25</points>
<connection>
<GID>198</GID>
<name>clock</name></connection>
<intersection>-30 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>35,-30,35,-25</points>
<connection>
<GID>194</GID>
<name>clock</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-5.5,67,-5.5</points>
<intersection>28 3</intersection>
<intersection>33.5 11</intersection>
<intersection>43 4</intersection>
<intersection>55 7</intersection>
<intersection>67 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-9.5,28,-5.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>43,-9.5,43,-5.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>55,-9.5,55,-5.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>67,-9.5,67,-5.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>33.5,-5.5,33.5,-3</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-22,35,-22</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<connection>
<GID>194</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-22,47,-22</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<connection>
<GID>196</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-22,59.5,-22</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<connection>
<GID>198</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,-22,71,-22</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<connection>
<GID>200</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-16,30.5,-15.5</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29,-15.5,30.5,-15.5</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-16,32.5,-15.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-15.5,33.5,-15.5</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-16,43.5,-15.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42,-15.5,43.5,-15.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-16,45.5,-15.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-15.5,46.5,-15.5</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-16,55.5,-15.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-15.5,55.5,-15.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-16,57.5,-15.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-15.5,58.5,-15.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-16,67.5,-15.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>66,-15.5,67.5,-15.5</points>
<connection>
<GID>217</GID>
<name>OUT</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-16,69.5,-15.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-15.5,70.5,-15.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-33.5,42,-22</points>
<connection>
<GID>223</GID>
<name>N_in3</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-22,42,-22</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>41 2</intersection>
<intersection>42 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>41,-22,41,-9.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-33.5,54,-22</points>
<connection>
<GID>225</GID>
<name>N_in3</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-22,54,-22</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection>
<intersection>54 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-22,53,-9.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-34,66,-22</points>
<connection>
<GID>227</GID>
<name>N_in3</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-22,66,-22</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>65.5 2</intersection>
<intersection>66 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>65.5,-22,65.5,-9.5</points>
<intersection>-22 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>65,-9.5,65.5,-9.5</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>65.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-34.5,79,-22</points>
<connection>
<GID>229</GID>
<name>N_in3</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-22,79,-22</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-9.5,47.5,-3</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-3,71.5,-3</points>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection>
<intersection>39 6</intersection>
<intersection>47.5 0</intersection>
<intersection>59.5 3</intersection>
<intersection>71.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59.5,-9.5,59.5,-3</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-3 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>71.5,-9.5,71.5,-3</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-3 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>39,-9.5,39,-3</points>
<intersection>-9.5 7</intersection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>34.5,-9.5,39,-9.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>39 6</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-9.5,30,-9.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-9.5,69.5,-9.5</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-9.5,32.5,-9.5</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<connection>
<GID>243</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-9.5,57.5,-9.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-9.5,45.5,-9.5</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<connection>
<GID>244</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>15.3,15.3856,269.515,-110.268</PageViewport>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>51,-2</position>
<gparam>LABEL_TEXT Universal Registor</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AE_DFF_LOW</type>
<position>34.5,-19.5</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>102 </output>
<input>
<ID>clock</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_DFF_LOW</type>
<position>49,-19.5</position>
<input>
<ID>IN_0</ID>107 </input>
<output>
<ID>OUT_0</ID>103 </output>
<input>
<ID>clock</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>255</ID>
<type>AE_DFF_LOW</type>
<position>65.5,-19.5</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>104 </output>
<input>
<ID>clock</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>256</ID>
<type>AE_DFF_LOW</type>
<position>82,-19.5</position>
<input>
<ID>IN_0</ID>109 </input>
<output>
<ID>OUT_0</ID>105 </output>
<input>
<ID>clock</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>258</ID>
<type>BB_CLOCK</type>
<position>25,-26.5</position>
<output>
<ID>CLK</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>260</ID>
<type>AE_MUX_4x1</type>
<position>35,-35</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>111 </input>
<input>
<ID>IN_3</ID>110 </input>
<output>
<ID>OUT</ID>106 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>98 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>261</ID>
<type>AE_MUX_4x1</type>
<position>49,-35</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_3</ID>112 </input>
<output>
<ID>OUT</ID>107 </output>
<input>
<ID>SEL_0</ID>95 </input>
<input>
<ID>SEL_1</ID>99 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_MUX_4x1</type>
<position>65,-35</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_3</ID>113 </input>
<output>
<ID>OUT</ID>108 </output>
<input>
<ID>SEL_0</ID>96 </input>
<input>
<ID>SEL_1</ID>100 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_MUX_4x1</type>
<position>82,-35</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_2</ID>115 </input>
<input>
<ID>IN_3</ID>114 </input>
<output>
<ID>OUT</ID>109 </output>
<input>
<ID>SEL_0</ID>97 </input>
<input>
<ID>SEL_1</ID>101 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_TOGGLE</type>
<position>17.5,-33</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_TOGGLE</type>
<position>17.5,-35.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>269</ID>
<type>GA_LED</type>
<position>35.5,-12.5</position>
<input>
<ID>N_in2</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>GA_LED</type>
<position>50,-12</position>
<input>
<ID>N_in2</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>GA_LED</type>
<position>66.5,-12</position>
<input>
<ID>N_in2</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>GA_LED</type>
<position>83,-12</position>
<input>
<ID>N_in2</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>DA_FROM</type>
<position>21.5,-33</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>279</ID>
<type>DA_FROM</type>
<position>21.5,-35.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>281</ID>
<type>DE_TO</type>
<position>28,-33</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>282</ID>
<type>DE_TO</type>
<position>42,-33</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>283</ID>
<type>DE_TO</type>
<position>58,-33</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>284</ID>
<type>DE_TO</type>
<position>74.5,-33</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s0</lparam></gate>
<gate>
<ID>285</ID>
<type>DE_TO</type>
<position>28,-35</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>286</ID>
<type>DE_TO</type>
<position>42,-35</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>287</ID>
<type>DE_TO</type>
<position>58,-35</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>288</ID>
<type>DE_TO</type>
<position>75,-35</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID s1</lparam></gate>
<gate>
<ID>290</ID>
<type>AA_TOGGLE</type>
<position>33,-46</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_TOGGLE</type>
<position>46.5,-46.5</position>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_TOGGLE</type>
<position>63,-46</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>293</ID>
<type>AA_TOGGLE</type>
<position>79.5,-46</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_TOGGLE</type>
<position>83.5,-46</position>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_TOGGLE</type>
<position>37,-46</position>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>30.5,-15</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID q1</lparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>45,-14.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID q2</lparam></gate>
<gate>
<ID>299</ID>
<type>DA_FROM</type>
<position>61.5,-14.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID q3</lparam></gate>
<gate>
<ID>300</ID>
<type>DA_FROM</type>
<position>78,-14.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID q4</lparam></gate>
<gate>
<ID>302</ID>
<type>DE_TO</type>
<position>85,-40.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID q4</lparam></gate>
<gate>
<ID>303</ID>
<type>DE_TO</type>
<position>68,-40</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID q3</lparam></gate>
<gate>
<ID>304</ID>
<type>DE_TO</type>
<position>52,-40</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID q2</lparam></gate>
<gate>
<ID>305</ID>
<type>DE_TO</type>
<position>38,-40</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID q1</lparam></gate>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-26.5,35.5,-22.5</points>
<connection>
<GID>253</GID>
<name>clock</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-26.5,83,-26.5</points>
<connection>
<GID>258</GID>
<name>CLK</name></connection>
<intersection>35.5 0</intersection>
<intersection>50 4</intersection>
<intersection>66.5 5</intersection>
<intersection>83 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83,-26.5,83,-22.5</points>
<connection>
<GID>256</GID>
<name>clock</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>50,-26.5,50,-22.5</points>
<connection>
<GID>254</GID>
<name>clock</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>66.5,-26.5,66.5,-22.5</points>
<connection>
<GID>255</GID>
<name>clock</name></connection>
<intersection>-26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>19.5,-33,19.5,-33</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<connection>
<GID>277</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>19.5,-35.5,19.5,-35.5</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-34,30,-33</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<connection>
<GID>260</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-34,44,-33</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<connection>
<GID>261</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-34,60,-33</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<connection>
<GID>262</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-34,77,-33</points>
<connection>
<GID>263</GID>
<name>SEL_0</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-33,77,-33</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-35,30,-35</points>
<connection>
<GID>260</GID>
<name>SEL_1</name></connection>
<connection>
<GID>285</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-35,44,-35</points>
<connection>
<GID>261</GID>
<name>SEL_1</name></connection>
<connection>
<GID>286</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-35,60,-35</points>
<connection>
<GID>262</GID>
<name>SEL_1</name></connection>
<connection>
<GID>287</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-35,77,-35</points>
<connection>
<GID>263</GID>
<name>SEL_1</name></connection>
<connection>
<GID>288</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-16.5,32.5,-15</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>35.5,-15,35.5,-13.5</points>
<connection>
<GID>269</GID>
<name>N_in2</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-15,35.5,-15</points>
<intersection>32.5 0</intersection>
<intersection>35.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-16.5,47,-14.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50,-14.5,50,-13</points>
<connection>
<GID>271</GID>
<name>N_in2</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,-14.5,50,-14.5</points>
<intersection>47 0</intersection>
<intersection>50 1</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-16.5,63.5,-14.5</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>66.5,-14.5,66.5,-13</points>
<connection>
<GID>273</GID>
<name>N_in2</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-14.5,66.5,-14.5</points>
<intersection>63.5 0</intersection>
<intersection>66.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-16.5,80,-14.5</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>83,-14.5,83,-13</points>
<connection>
<GID>275</GID>
<name>N_in2</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-14.5,83,-14.5</points>
<intersection>80 0</intersection>
<intersection>83 1</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-32,35,-27</points>
<connection>
<GID>260</GID>
<name>OUT</name></connection>
<intersection>-27 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32.5,-27,32.5,-22.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-27,35,-27</points>
<intersection>32.5 1</intersection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-32,49,-27</points>
<connection>
<GID>261</GID>
<name>OUT</name></connection>
<intersection>-27 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>47,-27,47,-22.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,-27,49,-27</points>
<intersection>47 1</intersection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-32,65,-27</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-27 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>63.5,-27,63.5,-22.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-27,65,-27</points>
<intersection>63.5 1</intersection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-32,82,-27</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>-27 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>80,-27,80,-22.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-27,82,-27</points>
<intersection>80 1</intersection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-41,32,-38</points>
<connection>
<GID>260</GID>
<name>IN_3</name></connection>
<intersection>-41 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>33,-44,33,-41</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,-41,33,-41</points>
<intersection>32 0</intersection>
<intersection>33 1</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-41,36,-38</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>-41 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>37,-44,37,-41</points>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36,-41,37,-41</points>
<intersection>36 0</intersection>
<intersection>37 1</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-41,46,-38</points>
<connection>
<GID>261</GID>
<name>IN_3</name></connection>
<intersection>-41 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46.5,-44.5,46.5,-41</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46,-41,46.5,-41</points>
<intersection>46 0</intersection>
<intersection>46.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-41,62,-38</points>
<connection>
<GID>262</GID>
<name>IN_3</name></connection>
<intersection>-41 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>63,-44,63,-41</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62,-41,63,-41</points>
<intersection>62 0</intersection>
<intersection>63 1</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-41,79,-38</points>
<connection>
<GID>263</GID>
<name>IN_3</name></connection>
<intersection>-41 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>79.5,-44,79.5,-41</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79,-41,79.5,-41</points>
<intersection>79 0</intersection>
<intersection>79.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-44,83.5,-41</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>81,-41,81,-38</points>
<connection>
<GID>263</GID>
<name>IN_2</name></connection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>81,-41,83.5,-41</points>
<intersection>81 1</intersection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-38.5,85,-38</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-38,68,-38</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<connection>
<GID>303</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-38,52,-38</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<connection>
<GID>304</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-38,38,-38</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<connection>
<GID>305</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 5>
<page 6>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 6>
<page 7>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 7>
<page 8>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 8>
<page 9>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 9></circuit>